// DESCRIPTION: Verilator: 
//
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2015 by Todd Strader.

interface foo_intf;
    logic a;
endinterface

function integer the_other_func (input integer val);
    return val;
endfunction

module t (/*AUTOARG*/);
   genvar the_genvar;
   generate
      for (the_genvar = 0; the_genvar < 4; the_genvar++) begin: foo_loop
         foo foo_inst();
      end
   endgenerate

   bar bar_inst();

   logic x;
   assign x = foo_loop[bar_inst.THE_LP].foo_inst.y;
endmodule

module foo();
    logic y;
endmodule

module bar();
    localparam THE_LP = 2;
endmodule

