// DESCRIPTION: Verilator: Verilog Test module
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2019 by Todd Strader.

`define CHECK(sig) \
        if (sig``_in != sig``_out) begin \
            $display(`"%%Error (%m) sig``_in (0x%0x) != sig``_out (0x%0x)`", \
                     sig``_in, sig``_out); \
            $stop; \
        end

module t (/*AUTOARG*/
   // Inputs
   clk
   );
   input clk;

    genvar x;
    generate
        for (x = 0; x < 2; x = x + 1) begin: gen_loop
            integer cyc = 0;
            logic [31:0] accum_in;
            logic [31:0] accum_out;
            logic accum_bypass;
            logic [31:0] accum_bypass_out;
            logic [31:0] accum_out_expect;
            logic [31:0] accum_bypass_out_expect;
            logic s1_in;
            logic s1_out;
            logic [1:0] s2_in;
            logic [1:0] s2_out;
            logic [7:0] s8_in;
            logic [7:0] s8_out;
            logic [32:0] s33_in;
            logic [32:0] s33_out;
            logic [63:0] s64_in;
            logic [63:0] s64_out;
            logic [64:0] s65_in;
            logic [64:0] s65_out;
            logic [128:0] s129_in;
            logic [128:0] s129_out;

            secret
            secret (
                .accum_in,
                .accum_out,
                .accum_bypass,
                .accum_bypass_out,
                .s1_in,
                .s1_out,
                .s2_in,
                .s2_out,
                .s8_in,
                .s8_out,
                .s33_in,
                .s33_out,
                .s64_in,
                .s64_out,
                .s65_in,
                .s65_out,
                .s129_in,
                .s129_out,
                .clk);

            always @(posedge clk) begin
`ifdef TEST_VERBOSE
                $display("[%0t] x=%0d, cyc=%0d accum_in=%0d accum_out=%0d accum_bypass_out=%0d",
                         $time, x, cyc, accum_in, accum_out, accum_bypass_out);
`endif
                cyc <= cyc + 1;
                accum_in <= accum_in + 5;
                accum_out_expect <= accum_in + accum_out_expect;
                if (cyc == 0) begin
                    accum_in <= x*100;
                    accum_bypass <= '0;
                end else if (cyc > 0) begin
                    if (accum_out_expect != accum_out) begin
                        $display("%%Error: (%m) accum_out expected %0d got %0d",
                                 accum_out_expect, accum_out);
                        $stop;
                    end
                    if (accum_bypass_out_expect != accum_bypass_out) begin
                        $display("%%Error: (%m) accum_bypass_out expected %0d got %0d",
                                 accum_bypass_out_expect, accum_bypass_out);
                        $stop;
                    end
                    `CHECK(s1)
                    `CHECK(s2)
                    `CHECK(s8)
                    `CHECK(s33)
                    `CHECK(s64)
                    `CHECK(s65)
                    `CHECK(s129)
                end

                if (cyc == 5) accum_bypass <= '1;

                if (cyc == 10) begin
                    $write("*-* All Finished *-*\n");
                    $finish;
                end
            end

            assign accum_bypass_out_expect = accum_bypass ? accum_in :
                                                accum_out_expect;
        end
    endgenerate

endmodule
